library verilog;
use verilog.vl_types.all;
entity lab_2_part1_vlg_sample_tst is
    port(
        Clk             : in     vl_logic;
        x               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab_2_part1_vlg_sample_tst;
