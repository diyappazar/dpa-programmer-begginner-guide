library verilog;
use verilog.vl_types.all;
entity lab_2_part2 is
    port(
        x               : in     vl_logic;
        Clk             : in     vl_logic;
        Y               : out    vl_logic
    );
end lab_2_part2;
