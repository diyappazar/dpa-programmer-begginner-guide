library verilog;
use verilog.vl_types.all;
entity lab_2_part2_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab_2_part2_vlg_check_tst;
